module lib

pub struct Enemy {
pub mut:
	dir Direction
	pos Pos
	value int
}
